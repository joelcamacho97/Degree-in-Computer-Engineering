`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:07:57 11/07/2018 
// Design Name: 
// Module Name:    Projeto2018 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Projeto2018(
    input EN,
    input I,
    output P,
    output G,
    output C
    );
	 
	 


endmodule
